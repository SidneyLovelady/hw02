magic
tech sky130A
magscale 1 2
timestamp 1680227980
<< nwell >>
rect 3020 1450 3530 1650
rect 5020 1450 5530 1650
rect 2080 980 6635 1450
<< pwell >>
rect 400 640 6160 920
rect 390 -280 6160 640
rect 390 -560 6150 -280
<< psubdiff >>
rect 510 -330 1910 -300
rect 510 -500 540 -330
rect 1880 -500 1910 -330
rect 510 -530 1910 -500
rect 3270 -370 4430 -300
rect 3270 -460 3340 -370
rect 4360 -460 4430 -370
rect 3270 -530 4430 -460
<< nsubdiff >>
rect 3110 1530 3460 1590
rect 3110 1420 3190 1530
rect 3380 1420 3460 1530
rect 3110 1360 3460 1420
rect 5070 1510 5480 1590
rect 5070 1410 5200 1510
rect 5360 1410 5480 1510
rect 5070 1340 5480 1410
<< psubdiffcont >>
rect 540 -500 1880 -330
rect 3340 -460 4360 -370
<< nsubdiffcont >>
rect 3190 1420 3380 1530
rect 5200 1410 5360 1510
<< locali >>
rect 5150 1510 5400 1540
rect 5150 1410 5200 1510
rect 5360 1410 5400 1510
rect 5150 1380 5400 1410
rect 510 -330 1910 -300
rect 510 -500 540 -330
rect 1880 -500 1910 -330
rect 510 -530 1910 -500
<< viali >>
rect 3170 1530 3400 1550
rect 3170 1420 3190 1530
rect 3190 1420 3380 1530
rect 3380 1420 3400 1530
rect 3170 1400 3400 1420
rect 540 -500 1880 -330
rect 3310 -370 4390 -340
rect 3310 -460 3340 -370
rect 3340 -460 4360 -370
rect 4360 -460 4390 -370
rect 3310 -490 4390 -460
<< metal1 >>
rect -302 1650 1158 1658
rect -302 1550 6448 1650
rect -302 1459 3170 1550
rect -302 1456 1158 1459
rect -302 1016 -44 1456
rect 2452 1320 2645 1459
rect 3020 1400 3170 1459
rect 3400 1459 6448 1550
rect 3400 1400 3530 1459
rect 2230 1106 2419 1235
rect 2454 1195 2643 1320
rect 3020 1310 3530 1400
rect 4161 1308 4354 1459
rect 5070 1340 5480 1459
rect 5579 1386 6440 1459
rect 5572 1341 6440 1386
rect 2841 1259 3987 1280
rect 2679 1244 3987 1259
rect 2456 1052 2645 1151
rect 2679 1115 4128 1244
rect 4163 1201 4352 1308
rect 2679 1070 3987 1115
rect 2679 1052 2877 1070
rect 4163 1060 4352 1161
rect 4392 1122 4581 1251
rect 5347 1232 5536 1233
rect 5012 1104 5536 1232
rect 5572 1187 6437 1341
rect -302 280 -23 1016
rect 2403 940 2877 1052
rect 4112 940 4404 1060
rect 5012 940 5413 1104
rect 5571 943 6436 1142
rect 6472 1101 6661 1230
rect 820 851 2877 940
rect 3300 912 5413 940
rect 591 649 780 778
rect 820 740 2800 851
rect 816 580 2796 696
rect 2839 651 2918 780
rect 3184 645 3266 774
rect 3300 740 5280 912
rect 3304 580 5284 691
rect 5328 653 5517 782
rect 816 496 5284 580
rect 5751 548 6144 943
rect 1475 491 5284 496
rect 1475 334 4633 491
rect 5425 480 5637 490
rect 5425 351 5719 480
rect 5752 441 5941 548
rect 1475 324 3510 334
rect -302 92 2120 280
rect -300 90 2120 92
rect 1888 74 2110 90
rect 1919 44 2110 74
rect 2463 47 3510 324
rect 1694 -126 1883 3
rect 1919 -40 2108 44
rect 2217 7 2382 8
rect 2143 -11 2382 7
rect 1917 -170 2106 -79
rect 2143 -122 2555 -11
rect 2587 -52 2979 47
rect 5425 5 5637 351
rect 5755 300 5944 397
rect 5977 356 6166 485
rect 3162 2 5637 5
rect 3162 -8 5644 2
rect 2217 -140 2555 -122
rect 1917 -208 2110 -170
rect 1920 -300 2110 -208
rect 2589 -217 2981 -96
rect 3016 -137 5644 -8
rect 3162 -153 5644 -137
rect 3162 -156 5461 -153
rect 2589 -219 2982 -217
rect 2590 -300 2982 -219
rect 5740 -300 5950 300
rect 510 -330 5950 -300
rect 510 -500 540 -330
rect 1880 -340 5950 -330
rect 1880 -490 3310 -340
rect 4390 -490 5950 -340
rect 1880 -500 5950 -490
rect 510 -530 5950 -500
use sky130_fd_pr__nfet_01v8_4W7PEP  sky130_fd_pr__nfet_01v8_4W7PEP_0
timestamp 1679528750
transform 0 1 5848 -1 0 417
box -73 -188 73 188
use sky130_fd_pr__nfet_01v8_UNLS5X  sky130_fd_pr__nfet_01v8_UNLS5X_0
timestamp 1679527038
transform 0 1 4297 -1 0 714
box -73 -1088 73 1088
use sky130_fd_pr__pfet_01v8_XGALHL  sky130_fd_pr__pfet_01v8_XGALHL_0
timestamp 1679526914
transform 0 1 4258 -1 0 1183
box -109 -200 109 200
use sky130_fd_pr__nfet_01v8_UNLS5X  XM1
timestamp 1679527038
transform 0 1 1810 -1 0 715
box -73 -1088 73 1088
use sky130_fd_pr__pfet_01v8_XGALHL  XM3
timestamp 1679526914
transform 0 1 2550 -1 0 1171
box -109 -200 109 200
use sky130_fd_pr__nfet_01v8_J2SMEF  XM5
timestamp 1679527038
transform 0 1 2784 -1 0 -75
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_4W7PEP  XM6
timestamp 1679528750
transform 0 1 2012 -1 0 -61
box -73 -188 73 188
use sky130_fd_pr__pfet_01v8_M6JSNY  XM8
timestamp 1679527038
transform 0 1 6003 -1 0 1163
box -109 -537 109 537
<< labels >>
rlabel metal1 -302 1456 1158 1658 1 VDD
port 1 n
rlabel metal1 591 649 780 778 1 Vinp
port 2 n
rlabel metal1 5328 653 5517 782 1 Vinn
port 3 n
rlabel metal1 2590 -530 2981 -96 1 VSS
port 4 n
rlabel metal1 5012 912 5413 1232 1 s1
port 5 n
rlabel metal1 5751 548 6144 1142 1 s2
port 6 n
<< end >>
