magic
tech sky130A
magscale 1 2
timestamp 1679530652
<< nwell >>
rect 2080 980 6635 1450
<< pwell >>
rect 400 -280 6160 920
<< metal1 >>
rect -302 1650 1158 1658
rect -302 1459 6448 1650
rect -302 1456 1158 1459
rect -302 1016 -44 1456
rect 2452 1320 2645 1459
rect 2230 1106 2419 1235
rect 2454 1195 2643 1320
rect 4161 1308 4354 1459
rect 5579 1386 6440 1459
rect 5572 1341 6440 1386
rect 2841 1259 3987 1280
rect 2679 1244 3987 1259
rect 2456 1052 2645 1151
rect 2679 1115 4128 1244
rect 4163 1201 4352 1308
rect 2679 1070 3987 1115
rect 2679 1052 2877 1070
rect 4163 1060 4352 1161
rect 4392 1122 4581 1251
rect 5347 1232 5536 1233
rect 5012 1104 5536 1232
rect 5572 1187 6437 1341
rect -302 272 -23 1016
rect 2403 940 2877 1052
rect 4112 940 4404 1060
rect 5012 940 5413 1104
rect 5571 943 6436 1142
rect 6472 1101 6661 1230
rect 820 851 2877 940
rect 3300 912 5413 940
rect 591 649 780 778
rect 820 740 2800 851
rect 816 580 2796 696
rect 2839 651 2918 780
rect 3184 645 3266 774
rect 3300 740 5280 912
rect 3304 580 5284 691
rect 5328 653 5517 782
rect 816 496 5284 580
rect 5751 548 6144 943
rect 1475 491 5284 496
rect 1475 334 4633 491
rect 5425 480 5637 490
rect 5425 351 5719 480
rect 5752 441 5941 548
rect 1475 324 3510 334
rect -302 251 1109 272
rect -302 198 2106 251
rect -302 105 2110 198
rect -302 92 1109 105
rect 1888 74 2110 105
rect 1919 44 2110 74
rect 2463 47 3510 324
rect 1694 -126 1883 3
rect 1919 -40 2108 44
rect 2217 7 2382 8
rect 2143 -11 2382 7
rect 1917 -208 2106 -79
rect 2143 -122 2555 -11
rect 2587 -52 2979 47
rect 5425 5 5637 351
rect 5755 268 5944 397
rect 5977 356 6166 485
rect 3162 2 5637 5
rect 3162 -8 5644 2
rect 2217 -140 2555 -122
rect 2589 -219 2981 -96
rect 3016 -137 5644 -8
rect 3162 -153 5644 -137
rect 3162 -156 5461 -153
use sky130_fd_pr__nfet_01v8_UNLS5X  XM1
timestamp 1679527038
transform 0 1 1810 -1 0 715
box -73 -1088 73 1088
use sky130_fd_pr__pfet_01v8_XGALHL  XM3
timestamp 1679526914
transform 0 1 2550 -1 0 1171
box -109 -200 109 200
use sky130_fd_pr__nfet_01v8_J2SMEF  XM5
timestamp 1679527038
transform 0 1 2784 -1 0 -75
box -73 -288 73 288
use sky130_fd_pr__nfet_01v8_4W7PEP  XM6
timestamp 1679528750
transform 0 1 2012 -1 0 -61
box -73 -188 73 188
use sky130_fd_pr__pfet_01v8_M6JSNY  XM8
timestamp 1679527038
transform 0 1 6003 -1 0 1163
box -109 -537 109 537
use sky130_fd_pr__nfet_01v8_4W7PEP  sky130_fd_pr__nfet_01v8_4W7PEP_0
timestamp 1679528750
transform 0 1 5848 -1 0 417
box -73 -188 73 188
use sky130_fd_pr__nfet_01v8_UNLS5X  sky130_fd_pr__nfet_01v8_UNLS5X_0
timestamp 1679527038
transform 0 1 4297 -1 0 714
box -73 -1088 73 1088
use sky130_fd_pr__pfet_01v8_XGALHL  sky130_fd_pr__pfet_01v8_XGALHL_0
timestamp 1679526914
transform 0 1 4258 -1 0 1183
box -109 -200 109 200
<< end >>
